`define addrWidth 8
`define dataWidth 8
